library verilog;
use verilog.vl_types.all;
entity Neander_vlg_vec_tst is
end Neander_vlg_vec_tst;
